module adc(
	input clk50,
	input [9:0]idata,
	output [39:0]odata,
	output wren
);

endmodule
