`ifndef DEF
`define DEF
typedef byte u8;
typedef int unsigned u32;
typedef logic [5:0]u6;
typedef logic [27:0]u28;
`endif
