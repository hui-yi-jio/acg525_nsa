`ifndef DEF
`define DEF
typedef byte u8;
typedef int unsigned u32;

`endif
