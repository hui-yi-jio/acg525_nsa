module rx(
	input rxclk, rxctl,
	input [3:0]rxd
);
	
endmodule
